// #############################################################################################################################
// VECTOR ALU
// 
// 向量计算时每个lane中一个
// #############################################################################################################################
module VECTOR_ALU#(parameter ADDR_WIDTH = 17,
                   parameter LEN = 32,
                   parameter BYTE_SIZE = 8,
                   parameter VECTOR_SIZE = 8,
                   parameter ENTRY_INDEX_SIZE = 3)
                  ();
    
endmodule
